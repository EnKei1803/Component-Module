/*
==================================================================================================
		 ____                      _    ____  _     _  __ _            
		| __ )  __ _ _ __ _ __ ___| |  / ___|| |__ (_)/ _| |_ ___ _ __ 
		|  _ \ / _` | '__| '__/ _ \ |  \___ \| '_ \| | |_| __/ _ \ '__|
		| |_) | (_| | |  | | |  __/ |   ___) | | | | |  _| ||  __/ |   
		|____/ \__,_|_|  |_|  \___|_|  |____/|_| |_|_|_|  \__\___|_|   
                                                                
==================================================================================================
*/
module shifter_32bits
(
	input logic		[31:0] A,		// Input
	input logic		[ 4:0] B,		// Shift n bits
	input logic		[ 1:0] Sel,		// Select mode Shift
	output logic	[31:0] Y			// Output 
);
/*
							|--------------------|-----------|--------------|
							|	 OPERATING MODE	|	 Left		|	Arithmetic	|
							|--------------------|-----------|--------------|
							|		SHIFT RIGHT		|		0		|		  0		|
							|--------------------|-----------|--------------|
							|			 ASR			|		0		|		  1		|
							|--------------------|-----------|--------------|
							|		SHIFT LEFT		|		1		|		  0		|
							|--------------------|-----------|--------------|
							|			 ASL			|		1		|		  1		|
							|--------------------|-----------|--------------|


*/

logic zero;
assign zero = 1'b0; 

logic [31:0] A1, A2, A3, A4, A5, A6;

// Data Reversal
MUX_2x1 MUX_2x1_DIR_1  (Sel[1], A[0],  A[31], A6[0]);
MUX_2x1 MUX_2x1_DIR_2  (Sel[1], A[1],  A[30], A6[1]);
MUX_2x1 MUX_2x1_DIR_3  (Sel[1], A[2],  A[29], A6[2]);
MUX_2x1 MUX_2x1_DIR_4  (Sel[1], A[3],  A[28], A6[3]);
MUX_2x1 MUX_2x1_DIR_5  (Sel[1], A[4],  A[27], A6[4]);
MUX_2x1 MUX_2x1_DIR_6  (Sel[1], A[5],  A[26], A6[5]);
MUX_2x1 MUX_2x1_DIR_7  (Sel[1], A[6],  A[25], A6[6]);
MUX_2x1 MUX_2x1_DIR_8  (Sel[1], A[7],  A[24], A6[7]);
MUX_2x1 MUX_2x1_DIR_9  (Sel[1], A[8],  A[23], A6[8]);
MUX_2x1 MUX_2x1_DIR_10 (Sel[1], A[9],  A[22], A6[9]);
MUX_2x1 MUX_2x1_DIR_11 (Sel[1], A[10], A[21], A6[10]);
MUX_2x1 MUX_2x1_DIR_12 (Sel[1], A[11], A[20], A6[11]);
MUX_2x1 MUX_2x1_DIR_13 (Sel[1], A[12], A[19], A6[12]);
MUX_2x1 MUX_2x1_DIR_14 (Sel[1], A[13], A[18], A6[13]);
MUX_2x1 MUX_2x1_DIR_15 (Sel[1], A[14], A[17], A6[14]);
MUX_2x1 MUX_2x1_DIR_16 (Sel[1], A[15], A[16], A6[15]);
MUX_2x1 MUX_2x1_DIR_17 (Sel[1], A[16], A[15], A6[16]);
MUX_2x1 MUX_2x1_DIR_18 (Sel[1], A[17], A[14], A6[17]);
MUX_2x1 MUX_2x1_DIR_19 (Sel[1], A[18], A[13], A6[18]);
MUX_2x1 MUX_2x1_DIR_20 (Sel[1], A[19], A[12], A6[19]);
MUX_2x1 MUX_2x1_DIR_21 (Sel[1], A[20], A[11], A6[20]);
MUX_2x1 MUX_2x1_DIR_22 (Sel[1], A[21], A[10], A6[21]);
MUX_2x1 MUX_2x1_DIR_23 (Sel[1], A[22], A[9],  A6[22]);
MUX_2x1 MUX_2x1_DIR_24 (Sel[1], A[23], A[8],  A6[23]);
MUX_2x1 MUX_2x1_DIR_25 (Sel[1], A[24], A[7],  A6[24]);
MUX_2x1 MUX_2x1_DIR_26 (Sel[1], A[25], A[6],  A6[25]);
MUX_2x1 MUX_2x1_DIR_27 (Sel[1], A[26], A[5],  A6[26]);
MUX_2x1 MUX_2x1_DIR_28 (Sel[1], A[27], A[4],  A6[27]);
MUX_2x1 MUX_2x1_DIR_29 (Sel[1], A[28], A[3],  A6[28]);
MUX_2x1 MUX_2x1_DIR_30 (Sel[1], A[29], A[2],  A6[29]);
MUX_2x1 MUX_2x1_DIR_31 (Sel[1], A[30], A[1],  A6[30]);
MUX_2x1 MUX_2x1_DIR_32 (Sel[1], A[31], A[0],  A6[31]);

// Select Arithmetic or Logical
// 1 : Arithmetic
// 0 : Logical

/*
					
										 0   A[31]
										_|____|_
							Sel[0]___\ 0  1 /
										 \____/
											 |
											AoL1	0
											_|____|_
								Sel[1]___\ 0  1 /
											 \____/
												|
											  AoL
									 _______________________
									|			|			|		|
									| Sel[1]	| Sel[0]	|  Y	|
									|________|________|_____|
									|			|			|		|
									| 	 0		|	 0		|  0	|
									|________|________|_____|		
									|			|			|		|
									| 	 0		| 	 1		|A[31]|
									|________|________|_____|	
									|			|			|		|
									| 	 1		|	 0		|  0	|
									|________|________|_____|		
									|			|			|		|
									| 	 1		| 	 1		|	0	|
									|________|________|_____|		
*/

logic AoL,AoL1;
MUX_2x1 MUX_2x1_AoL1 (Sel[0], zero, A[31], AoL1);
MUX_2x1 MUX_2x1_AoL  (Sel[1], AoL1, zero, AoL);

// B4 (16-bit shift)
MUX_2x1 MUX_2x1_1_1  (B[4], A6[0],  A6[16], A1[0]);
MUX_2x1 MUX_2x1_1_2  (B[4], A6[1],  A6[17], A1[1]);
MUX_2x1 MUX_2x1_1_3  (B[4], A6[2],  A6[18], A1[2]);
MUX_2x1 MUX_2x1_1_4  (B[4], A6[3],  A6[19], A1[3]);
MUX_2x1 MUX_2x1_1_5  (B[4], A6[4],  A6[20], A1[4]);
MUX_2x1 MUX_2x1_1_6  (B[4], A6[5],  A6[21], A1[5]);
MUX_2x1 MUX_2x1_1_7  (B[4], A6[6],  A6[22], A1[6]);
MUX_2x1 MUX_2x1_1_8  (B[4], A6[7],  A6[23], A1[7]);
MUX_2x1 MUX_2x1_1_9  (B[4], A6[8],  A6[24], A1[8]);
MUX_2x1 MUX_2x1_1_10 (B[4], A6[9],  A6[25], A1[9]);
MUX_2x1 MUX_2x1_1_11 (B[4], A6[10], A6[26], A1[10]);
MUX_2x1 MUX_2x1_1_12 (B[4], A6[11], A6[27], A1[11]);
MUX_2x1 MUX_2x1_1_13 (B[4], A6[12], A6[28], A1[12]);
MUX_2x1 MUX_2x1_1_14 (B[4], A6[13], A6[29], A1[13]);
MUX_2x1 MUX_2x1_1_15 (B[4], A6[14], A6[30], A1[14]);
MUX_2x1 MUX_2x1_1_16 (B[4], A6[15], A6[31], A1[15]);

MUX_2x1 MUX_2x1_1_17 (B[4], A6[16], AoL, A1[16]);
MUX_2x1 MUX_2x1_1_18 (B[4], A6[17], AoL, A1[17]);
MUX_2x1 MUX_2x1_1_19 (B[4], A6[18], AoL, A1[18]);
MUX_2x1 MUX_2x1_1_20 (B[4], A6[19], AoL, A1[19]);

MUX_2x1 MUX_2x1_1_21 (B[4], A6[20], AoL, A1[20]);
MUX_2x1 MUX_2x1_1_22 (B[4], A6[21], AoL, A1[21]);
MUX_2x1 MUX_2x1_1_23 (B[4], A6[22], AoL, A1[22]);
MUX_2x1 MUX_2x1_1_24 (B[4], A6[23], AoL, A1[23]);

MUX_2x1 MUX_2x1_1_25 (B[4], A6[24], AoL, A1[24]);
MUX_2x1 MUX_2x1_1_26 (B[4], A6[25], AoL, A1[25]);
MUX_2x1 MUX_2x1_1_27 (B[4], A6[26], AoL, A1[26]);
MUX_2x1 MUX_2x1_1_28 (B[4], A6[27], AoL, A1[27]);

MUX_2x1 MUX_2x1_1_29 (B[4], A6[28], AoL, A1[28]);
MUX_2x1 MUX_2x1_1_30 (B[4], A6[29], AoL, A1[29]);
MUX_2x1 MUX_2x1_1_31 (B[4], A6[30], AoL, A1[30]);
MUX_2x1 MUX_2x1_1_32 (B[4], A6[31], AoL, A1[31]);

// B3 (8-bit shift)
MUX_2x1 MUX_2x1_2_1  (B[3], A1[0],  A1[8],  A2[0]);
MUX_2x1 MUX_2x1_2_2  (B[3], A1[1],  A1[9],  A2[1]);
MUX_2x1 MUX_2x1_2_3  (B[3], A1[2],  A1[10], A2[2]);
MUX_2x1 MUX_2x1_2_4  (B[3], A1[3],  A1[11], A2[3]);
MUX_2x1 MUX_2x1_2_5  (B[3], A1[4],  A1[12], A2[4]);
MUX_2x1 MUX_2x1_2_6  (B[3], A1[5],  A1[13], A2[5]);
MUX_2x1 MUX_2x1_2_7  (B[3], A1[6],  A1[14], A2[6]);
MUX_2x1 MUX_2x1_2_8  (B[3], A1[7],  A1[15], A2[7]);
MUX_2x1 MUX_2x1_2_9  (B[3], A1[8],  A1[16], A2[8]);
MUX_2x1 MUX_2x1_2_10 (B[3], A1[9],  A1[17], A2[9]);
MUX_2x1 MUX_2x1_2_11 (B[3], A1[10], A1[18], A2[10]);
MUX_2x1 MUX_2x1_2_12 (B[3], A1[11], A1[19], A2[11]);
MUX_2x1 MUX_2x1_2_13 (B[3], A1[12], A1[20], A2[12]);
MUX_2x1 MUX_2x1_2_14 (B[3], A1[13], A1[21], A2[13]);
MUX_2x1 MUX_2x1_2_15 (B[3], A1[14], A1[22], A2[14]);
MUX_2x1 MUX_2x1_2_16 (B[3], A1[15], A1[23], A2[15]);
MUX_2x1 MUX_2x1_2_17 (B[3], A1[16], A1[24], A2[16]);
MUX_2x1 MUX_2x1_2_18 (B[3], A1[17], A1[25], A2[17]);
MUX_2x1 MUX_2x1_2_19 (B[3], A1[18], A1[26], A2[18]);
MUX_2x1 MUX_2x1_2_20 (B[3], A1[19], A1[27], A2[19]);
MUX_2x1 MUX_2x1_2_21 (B[3], A1[20], A1[28], A2[20]);
MUX_2x1 MUX_2x1_2_22 (B[3], A1[21], A1[29], A2[21]);
MUX_2x1 MUX_2x1_2_23 (B[3], A1[22], A1[30], A2[22]);
MUX_2x1 MUX_2x1_2_24 (B[3], A1[23], A1[31], A2[23]);

MUX_2x1 MUX_2x1_2_25 (B[3], A1[24], AoL, A2[24]);
MUX_2x1 MUX_2x1_2_26 (B[3], A1[25], AoL, A2[25]);
MUX_2x1 MUX_2x1_2_27 (B[3], A1[26], AoL, A2[26]);
MUX_2x1 MUX_2x1_2_28 (B[3], A1[27], AoL, A2[27]);

MUX_2x1 MUX_2x1_2_29 (B[3], A1[28], AoL, A2[28]);
MUX_2x1 MUX_2x1_2_30 (B[3], A1[29], AoL, A2[29]);
MUX_2x1 MUX_2x1_2_31 (B[3], A1[30], AoL, A2[30]);
MUX_2x1 MUX_2x1_2_32 (B[3], A1[31], AoL, A2[31]);

// B2 (4-bit shift)
MUX_2x1 MUX_2x1_3_1  (B[2], A2[0],  A2[4],  A3[0]);
MUX_2x1 MUX_2x1_3_2  (B[2], A2[1],  A2[5],  A3[1]);
MUX_2x1 MUX_2x1_3_3  (B[2], A2[2],  A2[6],  A3[2]);
MUX_2x1 MUX_2x1_3_4  (B[2], A2[3],  A2[7],  A3[3]);
MUX_2x1 MUX_2x1_3_5  (B[2], A2[4],  A2[8],  A3[4]);
MUX_2x1 MUX_2x1_3_6  (B[2], A2[5],  A2[9],  A3[5]);
MUX_2x1 MUX_2x1_3_7  (B[2], A2[6],  A2[10], A3[6]);
MUX_2x1 MUX_2x1_3_8  (B[2], A2[7],  A2[11], A3[7]);
MUX_2x1 MUX_2x1_3_9  (B[2], A2[8],  A2[12], A3[8]);
MUX_2x1 MUX_2x1_3_10 (B[2], A2[9],  A2[13], A3[9]);
MUX_2x1 MUX_2x1_3_11 (B[2], A2[10], A2[14], A3[10]);
MUX_2x1 MUX_2x1_3_12 (B[2], A2[11], A2[15], A3[11]);
MUX_2x1 MUX_2x1_3_13 (B[2], A2[12], A2[16], A3[12]);
MUX_2x1 MUX_2x1_3_14 (B[2], A2[13], A2[17], A3[13]);
MUX_2x1 MUX_2x1_3_15 (B[2], A2[14], A2[18], A3[14]);
MUX_2x1 MUX_2x1_3_16 (B[2], A2[15], A2[19], A3[15]);
MUX_2x1 MUX_2x1_3_17 (B[2], A2[16], A2[20], A3[16]);
MUX_2x1 MUX_2x1_3_18 (B[2], A2[17], A2[21], A3[17]);
MUX_2x1 MUX_2x1_3_19 (B[2], A2[18], A2[22], A3[18]);
MUX_2x1 MUX_2x1_3_20 (B[2], A2[19], A2[23], A3[19]);
MUX_2x1 MUX_2x1_3_21 (B[2], A2[20], A2[24], A3[20]);
MUX_2x1 MUX_2x1_3_22 (B[2], A2[21], A2[25], A3[21]);
MUX_2x1 MUX_2x1_3_23 (B[2], A2[22], A2[26], A3[22]);
MUX_2x1 MUX_2x1_3_24 (B[2], A2[23], A2[27], A3[23]);
MUX_2x1 MUX_2x1_3_25 (B[2], A2[24], A2[28], A3[24]);
MUX_2x1 MUX_2x1_3_26 (B[2], A2[25], A2[29], A3[25]);
MUX_2x1 MUX_2x1_3_27 (B[2], A2[26], A2[30], A3[26]);
MUX_2x1 MUX_2x1_3_28 (B[2], A2[27], A2[31], A3[27]);

MUX_2x1 MUX_2x1_3_29 (B[2], A2[28], AoL, A3[28]);
MUX_2x1 MUX_2x1_3_30 (B[2], A2[29], AoL, A3[29]);
MUX_2x1 MUX_2x1_3_31 (B[2], A2[30], AoL, A3[30]);
MUX_2x1 MUX_2x1_3_32 (B[2], A2[31], AoL, A3[31]);

// B1 (2-bit shift)
MUX_2x1 MUX_2x1_4_1  (B[1], A3[0],  A3[2],  A4[0]);
MUX_2x1 MUX_2x1_4_2  (B[1], A3[1],  A3[3],  A4[1]);
MUX_2x1 MUX_2x1_4_3  (B[1], A3[2],  A3[4],  A4[2]);
MUX_2x1 MUX_2x1_4_4  (B[1], A3[3],  A3[5],  A4[3]);
MUX_2x1 MUX_2x1_4_5  (B[1], A3[4],  A3[6],  A4[4]);
MUX_2x1 MUX_2x1_4_6  (B[1], A3[5],  A3[7],  A4[5]);
MUX_2x1 MUX_2x1_4_7  (B[1], A3[6],  A3[8],  A4[6]);
MUX_2x1 MUX_2x1_4_8  (B[1], A3[7],  A3[9],  A4[7]);
MUX_2x1 MUX_2x1_4_9  (B[1], A3[8],  A3[10], A4[8]);
MUX_2x1 MUX_2x1_4_10 (B[1], A3[9],  A3[11], A4[9]);
MUX_2x1 MUX_2x1_4_11 (B[1], A3[10], A3[12], A4[10]);
MUX_2x1 MUX_2x1_4_12 (B[1], A3[11], A3[13], A4[11]);
MUX_2x1 MUX_2x1_4_13 (B[1], A3[12], A3[14], A4[12]);
MUX_2x1 MUX_2x1_4_14 (B[1], A3[13], A3[15], A4[13]);
MUX_2x1 MUX_2x1_4_15 (B[1], A3[14], A3[16], A4[14]);
MUX_2x1 MUX_2x1_4_16 (B[1], A3[15], A3[17], A4[15]);
MUX_2x1 MUX_2x1_4_17 (B[1], A3[16], A3[18], A4[16]);
MUX_2x1 MUX_2x1_4_18 (B[1], A3[17], A3[19], A4[17]);
MUX_2x1 MUX_2x1_4_19 (B[1], A3[18], A3[20], A4[18]);
MUX_2x1 MUX_2x1_4_20 (B[1], A3[19], A3[21], A4[19]);
MUX_2x1 MUX_2x1_4_21 (B[1], A3[20], A3[22], A4[20]);
MUX_2x1 MUX_2x1_4_22 (B[1], A3[21], A3[23], A4[21]);
MUX_2x1 MUX_2x1_4_23 (B[1], A3[22], A3[24], A4[22]);
MUX_2x1 MUX_2x1_4_24 (B[1], A3[23], A3[25], A4[23]);
MUX_2x1 MUX_2x1_4_25 (B[1], A3[24], A3[26], A4[24]);
MUX_2x1 MUX_2x1_4_26 (B[1], A3[25], A3[27], A4[25]);
MUX_2x1 MUX_2x1_4_27 (B[1], A3[26], A3[28], A4[26]);
MUX_2x1 MUX_2x1_4_28 (B[1], A3[27], A3[29], A4[27]);
MUX_2x1 MUX_2x1_4_29 (B[1], A3[28], A3[30], A4[28]);
MUX_2x1 MUX_2x1_4_30 (B[1], A3[29], A3[31], A4[29]);

MUX_2x1 MUX_2x1_4_31 (B[1], A3[30], AoL, A4[30]);
MUX_2x1 MUX_2x1_4_32 (B[1], A3[31], AoL, A4[31]);

// B0 (1-bit shift)
MUX_2x1 MUX_2x1_5_1  (B[0], A4[0],  A4[1],  A5[0]);
MUX_2x1 MUX_2x1_5_2  (B[0], A4[1],  A4[2],  A5[1]);
MUX_2x1 MUX_2x1_5_3  (B[0], A4[2],  A4[3],  A5[2]);
MUX_2x1 MUX_2x1_5_4  (B[0], A4[3],  A4[4],  A5[3]);
MUX_2x1 MUX_2x1_5_5  (B[0], A4[4],  A4[5],  A5[4]);
MUX_2x1 MUX_2x1_5_6  (B[0], A4[5],  A4[6],  A5[5]);
MUX_2x1 MUX_2x1_5_7  (B[0], A4[6],  A4[7],  A5[6]);
MUX_2x1 MUX_2x1_5_8  (B[0], A4[7],  A4[8],  A5[7]);
MUX_2x1 MUX_2x1_5_9  (B[0], A4[8],  A4[9],  A5[8]);
MUX_2x1 MUX_2x1_5_10 (B[0], A4[9],  A4[10], A5[9]);
MUX_2x1 MUX_2x1_5_11 (B[0], A4[10], A4[11], A5[10]);
MUX_2x1 MUX_2x1_5_12 (B[0], A4[11], A4[12], A5[11]);
MUX_2x1 MUX_2x1_5_13 (B[0], A4[12], A4[13], A5[12]);
MUX_2x1 MUX_2x1_5_14 (B[0], A4[13], A4[14], A5[13]);
MUX_2x1 MUX_2x1_5_15 (B[0], A4[14], A4[15], A5[14]);
MUX_2x1 MUX_2x1_5_16 (B[0], A4[15], A4[16], A5[15]);
MUX_2x1 MUX_2x1_5_17 (B[0], A4[16], A4[17], A5[16]);
MUX_2x1 MUX_2x1_5_18 (B[0], A4[17], A4[18], A5[17]);
MUX_2x1 MUX_2x1_5_19 (B[0], A4[18], A4[19], A5[18]);
MUX_2x1 MUX_2x1_5_20 (B[0], A4[19], A4[20], A5[19]);
MUX_2x1 MUX_2x1_5_21 (B[0], A4[20], A4[21], A5[20]);
MUX_2x1 MUX_2x1_5_22 (B[0], A4[21], A4[22], A5[21]);
MUX_2x1 MUX_2x1_5_23 (B[0], A4[22], A4[23], A5[22]);
MUX_2x1 MUX_2x1_5_24 (B[0], A4[23], A4[24], A5[23]);
MUX_2x1 MUX_2x1_5_25 (B[0], A4[24], A4[25], A5[24]);
MUX_2x1 MUX_2x1_5_26 (B[0], A4[25], A4[26], A5[25]);
MUX_2x1 MUX_2x1_5_27 (B[0], A4[26], A4[27], A5[26]);
MUX_2x1 MUX_2x1_5_28 (B[0], A4[27], A4[28], A5[27]);
MUX_2x1 MUX_2x1_5_29 (B[0], A4[28], A4[29], A5[28]);
MUX_2x1 MUX_2x1_5_30 (B[0], A4[29], A4[30], A5[29]);
MUX_2x1 MUX_2x1_5_31 (B[0], A4[30], A4[31], A5[30]);

MUX_2x1 MUX_2x1_5_32 (B[0], A4[31], AoL, A5[31]);


// Data Reversal
MUX_2x1 MUX_2x1_OUT_1  (Sel[1], A5[0],  A5[31], Y[0]);
MUX_2x1 MUX_2x1_OUT_2  (Sel[1], A5[1],  A5[30], Y[1]);
MUX_2x1 MUX_2x1_OUT_3  (Sel[1], A5[2],  A5[29], Y[2]);
MUX_2x1 MUX_2x1_OUT_4  (Sel[1], A5[3],  A5[28], Y[3]);
MUX_2x1 MUX_2x1_OUT_5  (Sel[1], A5[4],  A5[27], Y[4]);
MUX_2x1 MUX_2x1_OUT_6  (Sel[1], A5[5],  A5[26], Y[5]);
MUX_2x1 MUX_2x1_OUT_7  (Sel[1], A5[6],  A5[25], Y[6]);
MUX_2x1 MUX_2x1_OUT_8  (Sel[1], A5[7],  A5[24], Y[7]);
MUX_2x1 MUX_2x1_OUT_9  (Sel[1], A5[8],  A5[23], Y[8]);
MUX_2x1 MUX_2x1_OUT_10 (Sel[1], A5[9],  A5[22], Y[9]);
MUX_2x1 MUX_2x1_OUT_11 (Sel[1], A5[10], A5[21], Y[10]);
MUX_2x1 MUX_2x1_OUT_12 (Sel[1], A5[11], A5[20], Y[11]);
MUX_2x1 MUX_2x1_OUT_13 (Sel[1], A5[12], A5[19], Y[12]);
MUX_2x1 MUX_2x1_OUT_14 (Sel[1], A5[13], A5[18], Y[13]);
MUX_2x1 MUX_2x1_OUT_15 (Sel[1], A5[14], A5[17], Y[14]);
MUX_2x1 MUX_2x1_OUT_16 (Sel[1], A5[15], A5[16], Y[15]);
MUX_2x1 MUX_2x1_OUT_17 (Sel[1], A5[16], A5[15], Y[16]);
MUX_2x1 MUX_2x1_OUT_18 (Sel[1], A5[17], A5[14], Y[17]);
MUX_2x1 MUX_2x1_OUT_19 (Sel[1], A5[18], A5[13], Y[18]);
MUX_2x1 MUX_2x1_OUT_20 (Sel[1], A5[19], A5[12], Y[19]);
MUX_2x1 MUX_2x1_OUT_21 (Sel[1], A5[20], A5[11], Y[20]);
MUX_2x1 MUX_2x1_OUT_22 (Sel[1], A5[21], A5[10], Y[21]);
MUX_2x1 MUX_2x1_OUT_23 (Sel[1], A5[22], A5[9],  Y[22]);
MUX_2x1 MUX_2x1_OUT_24 (Sel[1], A5[23], A5[8],  Y[23]);
MUX_2x1 MUX_2x1_OUT_25 (Sel[1], A5[24], A5[7],  Y[24]);
MUX_2x1 MUX_2x1_OUT_26 (Sel[1], A5[25], A5[6],  Y[25]);
MUX_2x1 MUX_2x1_OUT_27 (Sel[1], A5[26], A5[5],  Y[26]);
MUX_2x1 MUX_2x1_OUT_28 (Sel[1], A5[27], A5[4],  Y[27]);
MUX_2x1 MUX_2x1_OUT_29 (Sel[1], A5[28], A5[3],  Y[28]);
MUX_2x1 MUX_2x1_OUT_30 (Sel[1], A5[29], A5[2],  Y[29]);
MUX_2x1 MUX_2x1_OUT_31 (Sel[1], A5[30], A5[1],  Y[30]);
MUX_2x1 MUX_2x1_OUT_32 (Sel[1], A5[31], A5[0],  Y[31]);

endmodule 

