/*
==================================================================================================
           ___                                      ____           ___             
          |_ _|_ __   ___ _ __ ___  __ _ ___  ___  | __ ) _   _   / _ \ _ __   ___ 
           | || '_ \ / __| '__/ _ \/ _` / __|/ _ \ |  _ \| | | | | | | | '_ \ / _ \
           | || | | | (__| | |  __/ (_| \__ \  __/ | |_) | |_| | | |_| | | | |  __/
          |___|_| |_|\___|_|  \___|\__,_|___/\___| |____/ \__, |  \___/|_| |_|\___|
                                                          |___/                    
==================================================================================================
*/
module inc1
(
   input  logic [23:0] a,
   input  logic        cin,
   
   output logic [23:0] inc,
   output logic        cout 
   
);
logic [23:0] mask_string_s;

   string_gen  u_string_gen(
      .a    (a), 
      .cin  (cin), 
      .out  (mask_string_s), 
      .cout (cout)
   );

assign inc = mask_string_s ^ a;


endmodule

/*
==================================================================================================
        ____  _        _                ____                           _             
       / ___|| |_ _ __(_)_ __   __ _   / ___| ___ _ __   ___ _ __ __ _| |_ ___  _ __ 
       \___ \| __| '__| | '_ \ / _` | | |  _ / _ \ '_ \ / _ \ '__/ _` | __/ _ \| '__|
        ___) | |_| |  | | | | | (_| | | |_| |  __/ | | |  __/ | | (_| | || (_) | |   
       |____/ \__|_|  |_|_| |_|\__, |  \____|\___|_| |_|\___|_|  \__,_|\__\___/|_|   
                               |___/                                                 
==================================================================================================
*/

module string_gen
(
   input  logic [23:0] a,
   input  logic        cin,
   
   output logic [23:0] out,
   output logic        cout 
   
);

// ==================================================
//		            Extend size
// ==================================================

   logic [4:0] next_lsb;
   
   identical_block   u_out0   (.a(a[ 3: 0]),.lsb(cin),         .out(out[ 3: 0]), .next_lsb(next_lsb[0]) );   
   identical_block   u_out1   (.a(a[ 7: 4]),.lsb(next_lsb[0]), .out(out[ 7: 4]), .next_lsb(next_lsb[1]) );
   identical_block   u_out2   (.a(a[11: 8]),.lsb(next_lsb[1]), .out(out[11: 8]), .next_lsb(next_lsb[2]) );
   identical_block   u_out3   (.a(a[15:12]),.lsb(next_lsb[2]), .out(out[15:12]), .next_lsb(next_lsb[3]) );
   identical_block   u_out4   (.a(a[19:16]),.lsb(next_lsb[3]), .out(out[19:16]), .next_lsb(next_lsb[4]) );
   identical_block   u_out5   (.a(a[23:20]),.lsb(next_lsb[4]), .out(out[23:20]), .next_lsb(cout)        );


endmodule 

/*
==================================================================================================
              ___    _            _   _           _   ____  _            _    
             |_ _|__| | ___ _ __ | |_(_) ___ __ _| | | __ )| | ___   ___| | __
              | |/ _` |/ _ \ '_ \| __| |/ __/ _` | | |  _ \| |/ _ \ / __| |/ /
              | | (_| |  __/ | | | |_| | (_| (_| | | | |_) | | (_) | (__|   < 
             |___\__,_|\___|_| |_|\__|_|\___\__,_|_| |____/|_|\___/ \___|_|\_\
                                                                              
==================================================================================================
*/
module identical_block
(
   input  logic [3:0] a,
   input  logic       lsb,
   
   output logic [3:0] out,
   output logic       next_lsb 
   
);
   logic [3:0] pre_out;

   assign pre_out[0] = a[0];
   assign pre_out[1] = a[0] & a[1];
   assign pre_out[2] = a[0] & a[1] & a[2];
   assign pre_out[3] = a[0] & a[1] & a[2] & a[3];
   
// ==================================================
//		            Results
// ==================================================

   assign out[0]   = lsb;
   assign out[1]   = lsb & pre_out[0];
   assign out[2]   = lsb & pre_out[1];    
   assign out[3]   = lsb & pre_out[2]; 
   assign next_lsb = lsb & pre_out[3]; 

endmodule 